module res (
		output wire  ninit_done  // ninit_done.reset
	);
endmodule

