module rom (
		output wire [127:0] q,       //       q.dataout
		input  wire [7:0]   address, // address.address
		input  wire         clock    //   clock.clk
	);
endmodule

