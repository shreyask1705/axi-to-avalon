module vio (
		output wire [2:0] source,     //    sources.source
		input  wire       source_clk  // source_clk.clk
	);
endmodule

